package simPKG;


endpackage : simPKG
//  Package: sysPKG
//
package sysPKG;
    //  Group: Parameters
    parameter CLK_FREQ = 50_000_000;

    //  Group: Typedefs

endpackage: sysPKG
